class common;
	static mailbox gen2bfm=new();
	static virtual axi_interface vif;
	static string testname;
endclass

