`include "AXI_MASTER_interface.sv"
`include "AXI_common.sv"
`include "AXI_MASTER_tx.sv"
`include "AXI_MASTER_gen.sv"
`include "AXI_MASTER_bfm.sv"
`include "AXI_SLAVE_bfm.sv"
`include "AXI_MASTER_env.sv"
`include "AXI_MASTER_top.sv"

